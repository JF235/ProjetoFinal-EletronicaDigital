** Profile: "SCHEMATIC1-bias"  [ C:\Users\jfcmp\Documentos\Git\EE610 Projeto Final\parte04\flipflop-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../flipflop-pspicefiles/flipflop.lib" 
* From [PSPICE NETLIST] section of C:\Users\jfcmp\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 50ns 0 5p 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
