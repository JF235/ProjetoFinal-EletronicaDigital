** Profile: "SCHEMATIC1-inversor"  [ C:\Users\jfcmp\Documentos\Git\EE610 Projeto Final\parte01\ee610_projeto_final-PSpiceFiles\SCHEMATIC1\inversor.sim ] 

** Creating circuit file "inversor.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ee610_projeto_final-pspicefiles/ee610_projeto_final.lib" 
.LIB "../../../ee610_projeto_final-pspicefiles/pinv.lib" 
.LIB "../../../ee610_projeto_final-pspicefiles/ninv.lib" 
* From [PSPICE NETLIST] section of C:\Users\jfcmp\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VI 0 3 0.001 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
