** Profile: "OSCILADOR-bias"  [ c:\users\jfcmp\documentos\git\ee610 projeto final\parte03\oscilador-pspicefiles\oscilador\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../oscilador-pspicefiles/oscilador.lib" 
* From [PSPICE NETLIST] section of C:\Users\jfcmp\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 20ns 0 1ps 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\OSCILADOR.net" 


.END
