** Profile: "Latch-Latch"  [ c:\users\jfcmp\documentos\git\ee610 projeto final\parte01\ee610_projeto_final-PSpiceFiles\Latch\Latch.sim ] 

** Creating circuit file "Latch.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ee610_projeto_final-pspicefiles/ee610_projeto_final.lib" 
.LIB "../../../ee610_projeto_final-pspicefiles/pinv.lib" 
.LIB "../../../ee610_projeto_final-pspicefiles/ninv.lib" 
* From [PSPICE NETLIST] section of C:\Users\jfcmp\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2ns 0 0.004ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Latch.net" 


.END
